module deneme_03(in,in1,outp);
input in,in1;
output outp;
assign outp=in & in1;
endmodule
