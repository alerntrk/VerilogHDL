module andGate(out,in,in1);
input in,in1;
output out;
assign out=in&in1;
endmodule
