module notGate(in,outp);
	input in;
	output outp;
	assign outp=~in;
endmodule
